module mojo_top(
    // 50MHz clock input
    input clk,
    // Input from reset button (active low)
    input rst_n,
    // cclk input from AVR, high when AVR is ready
    input cclk,
    // Outputs to the 8 onboard LEDs
    output[7:0]led,
    // AVR SPI connections
    output spi_miso,
    input spi_ss,
    input spi_mosi,
    input spi_sck,
    // AVR ADC channel select
    output [3:0] spi_channel,
    // Serial connections
    input avr_tx, // AVR Tx => FPGA Rx
    output avr_rx, // AVR Rx => FPGA Tx
    input avr_rx_busy, // AVR Rx buffer full
	 //addeed output for external interface with servo
	 output servo
    );

wire rst = ~rst_n; // make reset active high

// these signals should be high-z when not used
assign spi_miso = 1'bz; 
assign avr_rx = 1'bz; 
assign spi_channel = 4'bzzzz;

 assign led = 8'b0;// sending zeros to the leds
   
 wire [7:0] servo_position; //creating a 8 bit controller for 256 positions in the servomotor
   
	//instantiated counter and servocontroller
  counter #(.CTR_LEN(28)) servoCounter (
    .clk(clk),
    .rst(rst),
    .value(servo_position)
  );
   
  servo myServoController (
    .clk(clk),
    .rst(rst),
    .position(servo_position),
    .servo(servo)
  );
  
endmodule 
